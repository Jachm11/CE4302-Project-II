module RAM_1p_8g_20a_128b
(
	input logic [19:0] address, // 20 bits de direccion => 16 bits para las sub RAMs y 4 bits para tener 16 sub RAMs
	input logic [127:0] data_in,
	input logic [15:0] byte_enablers,
	
	input logic write_enable,
	input logic clock,
	
	output logic [127:0] data_out
);
	logic [3:0] offset;
	logic [15:0] address_without_offset;
	assign {address_without_offset, offset} = address;

	logic [15:0][15:0] sub_addresses;
	Address_offset_16_byte AO
	(
		.address_without_offset(address_without_offset),
		.offset(offset),

		.sub_address_0(sub_addresses[0]),
		.sub_address_1(sub_addresses[1]),
		.sub_address_2(sub_addresses[2]),
		.sub_address_3(sub_addresses[3]),
		.sub_address_4(sub_addresses[4]),
		.sub_address_5(sub_addresses[5]),
		.sub_address_6(sub_addresses[6]),
		.sub_address_7(sub_addresses[7]),
		.sub_address_8(sub_addresses[8]),
		.sub_address_9(sub_addresses[9]),
		.sub_address_10(sub_addresses[10]),
		.sub_address_11(sub_addresses[11]),
		.sub_address_12(sub_addresses[12]),
		.sub_address_13(sub_addresses[13]),
		.sub_address_14(sub_addresses[14]),
		.sub_address_15(sub_addresses[15])
	);
	
	logic [127:0] shifted_data_in;
	Circular_shifter_left_byte_N #(.N(128)) cslb
	(
		.shifting(data_in),
		.shift_amount(offset),

		.shifted(shifted_data_in)
	);
	
	logic [15:0] shifted_byte_enablers;
	assign shifted_byte_enablers = (write_enable) ? (byte_enablers << offset) : 16'b0;

	logic [127:0] data_out_aux;
	
	// Sub RAMs
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_0	
	(
		.address(sub_addresses[0]),
		.clock(clock),
		.data(shifted_data_in[7:0]),
		.wren(shifted_byte_enablers[0]),

		.q(data_out_aux[7:0])
	);
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_1
	(
		.address(sub_addresses[1]),
		.clock(clock),
		.data(shifted_data_in[15:8]),
		.wren(shifted_byte_enablers[1]),

		.q(data_out_aux[15:8])
	);
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_2
	(
		.address(sub_addresses[2]),
		.clock(clock),
		.data(shifted_data_in[23:16]),
		.wren(shifted_byte_enablers[2]),

		.q(data_out_aux[23:16])
	);
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_3
	(
		.address(sub_addresses[3]),
		.clock(clock),
		.data(shifted_data_in[31:24]),
		.wren(shifted_byte_enablers[3]),

		.q(data_out_aux[31:24])
	);
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_4
	(
		.address(sub_addresses[4]),
		.clock(clock),
		.data(shifted_data_in[39:32]),
		.wren(shifted_byte_enablers[4]),

		.q(data_out_aux[39:32])
	);
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_5
	(
		.address(sub_addresses[5]),
		.clock(clock),
		.data(shifted_data_in[47:40]),
		.wren(shifted_byte_enablers[5]),

		.q(data_out_aux[47:40])
	);
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_6
	(
		.address(sub_addresses[6]),
		.clock(clock),
		.data(shifted_data_in[55:48]),
		.wren(shifted_byte_enablers[6]),

		.q(data_out_aux[55:48])
	);
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_7
	(
		.address(sub_addresses[7]),
		.clock(clock),
		.data(shifted_data_in[63:56]),
		.wren(shifted_byte_enablers[7]),

		.q(data_out_aux[63:56])
	);
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_8
	(
		.address(sub_addresses[8]),
		.clock(clock),
		.data(shifted_data_in[71:64]),
		.wren(shifted_byte_enablers[8]),

		.q(data_out_aux[71:64])
	);
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_9
	(
		.address(sub_addresses[9]),
		.clock(clock),
		.data(shifted_data_in[79:72]),
		.wren(shifted_byte_enablers[9]),

		.q(data_out_aux[79:72])
	);
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_10
	(
		.address(sub_addresses[10]),
		.clock(clock),
		.data(shifted_data_in[87:80]),
		.wren(shifted_byte_enablers[10]),

		.q(data_out_aux[87:80])
	);
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_11
	(
		.address(sub_addresses[11]),
		.clock(clock),
		.data(shifted_data_in[95:88]),
		.wren(shifted_byte_enablers[11]),

		.q(data_out_aux[95:88])
	);
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_12
	(
		.address(sub_addresses[12]),
		.clock(clock),
		.data(shifted_data_in[103:96]),
		.wren(shifted_byte_enablers[12]),

		.q(data_out_aux[103:96])
	);
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_13
	(
		.address(sub_addresses[13]),
		.clock(clock),
		.data(shifted_data_in[111:104]),
		.wren(shifted_byte_enablers[13]),

		.q(data_out_aux[111:104])
	);
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_14
	(
		.address(sub_addresses[14]),
		.clock(clock),
		.data(shifted_data_in[119:112]),
		.wren(shifted_byte_enablers[14]),

		.q(data_out_aux[119:112])
	);
	RAM_1p_8w_16a_8b_from_file #(.PATH("/home/jachm/Documents/Repos/CE4302-Project-II/cpu+hdmi/src/Memory/Mifs/data_null/16a_8g_empty_init_file.mif")) sub_RAM_15
	(
		.address(sub_addresses[15]),
		.clock(clock),
		.data(shifted_data_in[127:120]),
		.wren(shifted_byte_enablers[15]),

		.q(data_out_aux[127:120])
	);

	Circular_shifter_right_byte_N #(.N(128)) csrb
	(
		.shifting(data_out_aux),
		.shift_amount(offset),

		.shifted(data_out)
	);
endmodule
/*
RAM_1p_8g_20a_128b RAM
(
	.address(),
	.data_in(),
	.byte_enablers(),
	.write_enable(),

	.clock(),

	.data_out()
);
*/